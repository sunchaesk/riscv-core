`timescale 1ns / 1ps

module alu_tb;
   // declare inputs
   reg [31:0] in_a, in_b;
   reg [3:0]  alu_control;

   // declare outputs
   reg [31:0] alu_result;
   reg        zero_flag;


endmodule
